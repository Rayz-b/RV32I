module adder(output  [31:0] y,input   [31:0] a, b);
     assign y = a + b;
endmodule